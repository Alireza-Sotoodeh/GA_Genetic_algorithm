$date
   Wed Aug 20 20:44:49 2025
$end
$version
  2019.2
$end
$timescale
  1ps
$end
$scope module lsfr_random_TB $end
$var reg 1 ! CLK_generator $end
$var reg 1 " RST $end
$var reg 32 # error_count $end
$var reg 32 $ test_count $end
$scope module intf $end
$var wire 1 % clk $end
$var wire 1 & rst $end
$var reg 1 ' start_lfsr $end
$var reg 58 ( seed_in [57:0] $end
$var reg 1 ) load_seed $end
$var reg 16 * random_out [15:0] $end
$upscope $end
$scope module DUT $end
$var wire 1 + clk $end
$var wire 1 , rst_n $end
$var wire 1 - start_lfsr $end
$var wire 58 . seed_in [57:0] $end
$var wire 1 / load_seed $end
$var reg 16 0 random_out [15:0] $end
$var reg 16 1 lfsr1 [15:0] $end
$var reg 15 2 lfsr2 [14:0] $end
$var reg 14 3 lfsr3 [13:0] $end
$var reg 13 4 lfsr4 [12:0] $end
$var reg 1 5 fb1 $end
$var reg 1 6 fb2 $end
$var reg 1 7 fb3 $end
$var reg 1 8 fb4 $end
$var reg 16 9 combined [15:0] $end
$var parameter 32 : WIDTH1 [31:0] $end
$var parameter 32 ; WIDTH2 [31:0] $end
$var parameter 32 < WIDTH3 [31:0] $end
$var parameter 32 = WIDTH4 [31:0] $end
$var parameter 16 > defualtSeed1 [15:0] $end
$var parameter 15 ? defualtSeed2 [14:0] $end
$var parameter 14 @ defualtSeed3 [13:0] $end
$var parameter 13 A defualtSeed4 [12:0] $end
$upscope $end
$scope task generator $end
$var reg 32 B num_tests $end
$scope begin Block77_3 $end
$var reg 32 C i $end
$upscope $end
$upscope $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0!
0"
b0 #
b0 $
0%
0&
x'
bx (
x)
bx *
0+
1,
x-
bx .
x/
bx 0
bx 1
bx 2
bx 3
bx 4
x5
x6
x7
x8
bx 9
b10000 :
b1111 ;
b1110 <
b1101 =
b1010110011100001 >
b11101111101110 ?
b10101110101101 @
b1110110101101 A
b0 B
b0 C
$end
#1000
1!
1%
1+
#2000
0!
0%
0+
#3000
1!
1%
1+
#4000
0!
1"
0%
1&
b1010100000110101 *
0+
0,
b1010100000110101 0
b1010110011100001 1
b11101111101110 2
b10101110101101 3
b1110110101101 4
15
06
07
18
b1010000100001111 9
#5000
1!
1%
1+
#6000
0!
0%
0+
#7000
1!
1%
1+
#8000
0!
0%
0+
#9000
1!
1%
1+
#10000
0!
0%
0+
#11000
1!
1%
1+
#12000
0!
0%
0+
#13000
1!
1%
1+
#14000
0!
0%
0+
#15000
1!
1%
1+
#16000
0!
0%
0+
#17000
1!
1%
1+
#18000
0!
0%
0+
#19000
1!
1%
1+
#20000
0!
0%
0+
#21000
1!
1%
1+
#22000
0!
0%
0+
#23000
1!
1%
1+
#24000
0!
0%
0+
#25000
1!
1%
1+
#26000
0!
0%
0+
#27000
1!
1%
1+
#28000
0!
0%
0+
#29000
1!
1%
1+
#30000
0!
0%
0+
#31000
1!
1%
1+
#32000
0!
0%
0+
#33000
1!
1%
1+
#34000
0!
0%
0+
#35000
1!
1%
1+
#36000
0!
0%
0+
#37000
1!
1%
1+
#38000
0!
0%
0+
#39000
1!
1%
1+
#40000
0!
0%
0+
#41000
1!
1%
1+
#42000
0!
0%
0+
#43000
1!
1%
1+
#44000
0!
0%
0+
#45000
1!
1%
1+
#46000
0!
0%
0+
#47000
1!
1%
1+
#48000
0!
0%
0+
#49000
1!
1%
1+
#50000
0!
0%
0+
#51000
1!
1%
1+
#52000
0!
0%
0+
#53000
1!
1%
1+
#54000
0!
0%
0+
#55000
1!
1%
1+
#56000
0!
0%
0+
#57000
1!
1%
1+
#58000
0!
0%
0+
#59000
1!
1%
1+
#60000
0!
0%
0+
#61000
1!
1%
1+
#62000
0!
0%
0+
#63000
1!
1%
1+
#64000
0!
0%
0+
#65000
1!
1%
1+
#66000
0!
0%
0+
#67000
1!
1%
1+
#68000
0!
0%
0+
#69000
1!
1%
1+
#70000
0!
0%
0+
#71000
1!
1%
1+
#72000
0!
0%
0+
#73000
1!
1%
1+
#74000
0!
0%
0+
#75000
1!
1%
1+
#76000
0!
0%
0+
#77000
1!
1%
1+
#78000
0!
0%
0+
#79000
1!
1%
1+
#80000
0!
0%
0+
#81000
1!
1%
1+
#82000
0!
0%
0+
#83000
1!
1%
1+
#84000
0!
0%
0+
#85000
1!
1%
1+
#86000
0!
0%
0+
#87000
1!
1%
1+
#88000
0!
0%
0+
#89000
1!
1%
1+
#90000
0!
0%
0+
#91000
1!
1%
1+
#92000
0!
0%
0+
#93000
1!
1%
1+
#94000
0!
0%
0+
#95000
1!
1%
1+
#96000
0!
0%
0+
#97000
1!
1%
1+
#98000
0!
0%
0+
#99000
1!
1%
1+
#100000
0!
0%
0+
#101000
1!
1%
1+
#102000
0!
0%
0+
#103000
1!
1%
1+
#104000
0!
0%
0+
#105000
1!
1%
1+
#106000
0!
0%
0+
#107000
1!
1%
1+
#108000
0!
0%
0+
#109000
1!
1%
1+
#110000
0!
0%
0+
#111000
1!
1%
1+
#112000
0!
0%
0+
#113000
1!
1%
1+
#114000
0!
0%
0+
#115000
1!
1%
1+
#116000
0!
0%
0+
#117000
1!
1%
1+
#118000
0!
0%
0+
#119000
1!
1%
1+
#120000
0!
0%
0+
#121000
1!
1%
1+
#122000
0!
0%
0+
#123000
1!
1%
1+
#124000
0!
0%
0+
#125000
1!
1%
1+
#126000
0!
0%
0+
#127000
1!
1%
1+
#128000
0!
0%
0+
#129000
1!
1%
1+
#130000
0!
0%
0+
#131000
1!
1%
1+
#132000
0!
0%
0+
#133000
1!
1%
1+
#134000
0!
0%
0+
#135000
1!
1%
1+
#136000
0!
0%
0+
#137000
1!
1%
1+
#138000
0!
0%
0+
#139000
1!
1%
1+
#140000
0!
0%
0+
#141000
1!
1%
1+
#142000
0!
0%
0+
#143000
1!
1%
1+
#144000
0!
0%
0+
#145000
1!
1%
1+
#146000
0!
0%
0+
#147000
1!
1%
1+
#148000
0!
0%
0+
#149000
1!
1%
1+
#150000
0!
0%
0+
#151000
1!
1%
1+
#152000
0!
0%
0+
#153000
1!
1%
1+
#154000
0!
0%
0+
#155000
1!
1%
1+
#156000
0!
0%
0+
#157000
1!
1%
1+
#158000
0!
0%
0+
#159000
1!
1%
1+
#160000
0!
0%
0+
#161000
1!
1%
1+
#162000
0!
0%
0+
#163000
1!
1%
1+
#164000
0!
0%
0+
#165000
1!
1%
1+
#166000
0!
0%
0+
#167000
1!
1%
1+
#168000
0!
0%
0+
#169000
1!
1%
1+
#170000
0!
0%
0+
#171000
1!
1%
1+
#172000
0!
0%
0+
#173000
1!
1%
1+
#174000
0!
0%
0+
#175000
1!
1%
1+
#176000
0!
0%
0+
#177000
1!
1%
1+
#178000
0!
0%
0+
#179000
1!
1%
1+
#180000
0!
0%
0+
#181000
1!
1%
1+
#182000
0!
0%
0+
#183000
1!
1%
1+
#184000
0!
0%
0+
#185000
1!
1%
1+
#186000
0!
0%
0+
#187000
1!
1%
1+
#188000
0!
0%
0+
#189000
1!
1%
1+
#190000
0!
0%
0+
#191000
1!
1%
1+
#192000
0!
0%
0+
#193000
1!
1%
1+
#194000
0!
0%
0+
#195000
1!
1%
1+
#196000
0!
0%
0+
#197000
1!
1%
1+
#198000
0!
0%
0+
#199000
1!
1%
1+
#200000
0!
0%
0+
#201000
1!
1%
1+
#202000
0!
0%
0+
#203000
1!
1%
1+
#204000
0!
0%
0+
#205000
1!
1%
1+
#206000
0!
0%
0+
#207000
1!
1%
1+
#208000
0!
0%
0+
#209000
1!
1%
1+
#210000
0!
0%
0+
#211000
1!
1%
1+
#212000
0!
0%
0+
#213000
1!
1%
1+
#214000
0!
0%
0+
#215000
1!
1%
1+
#216000
0!
0%
0+
#217000
1!
1%
1+
#218000
0!
0%
0+
#219000
1!
1%
1+
#220000
0!
0%
0+
#221000
1!
1%
1+
#222000
0!
0%
0+
#223000
1!
1%
1+
#224000
0!
0%
0+
#225000
1!
1%
1+
#226000
0!
0%
0+
#227000
1!
1%
1+
#228000
0!
0%
0+
#229000
1!
1%
1+
#230000
0!
0%
0+
#231000
1!
1%
1+
#232000
0!
0%
0+
#233000
1!
1%
1+
#234000
0!
0%
0+
#235000
1!
1%
1+
#236000
0!
0%
0+
#237000
1!
1%
1+
#238000
0!
0%
0+
#239000
1!
1%
1+
#240000
0!
0%
0+
#241000
1!
1%
1+
#242000
0!
0%
0+
#243000
1!
1%
1+
#244000
0!
0%
0+
#245000
1!
1%
1+
#246000
0!
0%
0+
#247000
1!
1%
1+
#248000
0!
0%
0+
#249000
1!
1%
1+
#250000
0!
0%
0+
#251000
1!
1%
1+
#252000
0!
0%
0+
#253000
1!
1%
1+
#254000
0!
0%
0+
#255000
1!
1%
1+
#256000
0!
0%
0+
#257000
1!
1%
1+
#258000
0!
0%
0+
#259000
1!
1%
1+
#260000
0!
0%
0+
#261000
1!
1%
1+
#262000
0!
0%
0+
#263000
1!
1%
1+
#264000
0!
0%
0+
#265000
1!
1%
1+
#266000
0!
0%
0+
#267000
1!
1%
1+
#268000
0!
0%
0+
#269000
1!
1%
1+
#270000
0!
0%
0+
#271000
1!
1%
1+
#272000
0!
0%
0+
#273000
1!
1%
1+
#274000
0!
0%
0+
#275000
1!
1%
1+
#276000
0!
0%
0+
#277000
1!
1%
1+
#278000
0!
0%
0+
#279000
1!
1%
1+
#280000
0!
0%
0+
#281000
1!
1%
1+
#282000
0!
0%
0+
#283000
1!
1%
1+
#284000
0!
0%
0+
#285000
1!
1%
1+
#286000
0!
0%
0+
#287000
1!
1%
1+
#288000
0!
0%
0+
#289000
1!
1%
1+
#290000
0!
0%
0+
#291000
1!
1%
1+
#292000
0!
0%
0+
#293000
1!
1%
1+
#294000
0!
0%
0+
#295000
1!
1%
1+
#296000
0!
0%
0+
#297000
1!
1%
1+
#298000
0!
0%
0+
#299000
1!
1%
1+
#300000
0!
0%
0+
#301000
1!
1%
1+
#302000
0!
0%
0+
#303000
1!
1%
1+
#304000
0!
0%
0+
#305000
1!
1%
1+
#306000
0!
0%
0+
#307000
1!
1%
1+
#308000
0!
0%
0+
#309000
1!
1%
1+
#310000
0!
0%
0+
#311000
1!
1%
1+
#312000
0!
0%
0+
#313000
1!
1%
1+
#314000
0!
0%
0+
#315000
1!
1%
1+
#316000
0!
0%
0+
#317000
1!
1%
1+
#318000
0!
0%
0+
#319000
1!
1%
1+
#320000
0!
0%
0+
#321000
1!
1%
1+
#322000
0!
0%
0+
#323000
1!
1%
1+
#324000
0!
0%
0+
#325000
1!
1%
1+
#326000
0!
0%
0+
#327000
1!
1%
1+
#328000
0!
0%
0+
#329000
1!
1%
1+
#330000
0!
0%
0+
#331000
1!
1%
1+
#332000
0!
0%
0+
#333000
1!
1%
1+
#334000
0!
0%
0+
#335000
1!
1%
1+
#336000
0!
0%
0+
#337000
1!
1%
1+
#338000
0!
0%
0+
#339000
1!
1%
1+
#340000
0!
0%
0+
#341000
1!
1%
1+
#342000
0!
0%
0+
#343000
1!
1%
1+
#344000
0!
0%
0+
#345000
1!
1%
1+
#346000
0!
0%
0+
#347000
1!
1%
1+
#348000
0!
0%
0+
#349000
1!
1%
1+
#350000
0!
0%
0+
#351000
1!
1%
1+
#352000
0!
0%
0+
#353000
1!
1%
1+
#354000
0!
0%
0+
#355000
1!
1%
1+
#356000
0!
0%
0+
#357000
1!
1%
1+
#358000
0!
0%
0+
#359000
1!
1%
1+
#360000
0!
0%
0+
#361000
1!
1%
1+
#362000
0!
0%
0+
#363000
1!
1%
1+
#364000
0!
0%
0+
#365000
1!
1%
1+
#366000
0!
0%
0+
#367000
1!
1%
1+
#368000
0!
0%
0+
#369000
1!
1%
1+
#370000
0!
0%
0+
#371000
1!
1%
1+
#372000
0!
0%
0+
#373000
1!
1%
1+
#374000
0!
0%
0+
#375000
1!
1%
1+
#376000
0!
0%
0+
#377000
1!
1%
1+
#378000
0!
0%
0+
#379000
1!
1%
1+
#380000
0!
0%
0+
#381000
1!
1%
1+
#382000
0!
0%
0+
#383000
1!
1%
1+
#384000
0!
0%
0+
#385000
1!
1%
1+
#386000
0!
0%
0+
#387000
1!
1%
1+
#388000
0!
0%
0+
#389000
1!
1%
1+
#390000
0!
0%
0+
#391000
1!
1%
1+
#392000
0!
0%
0+
#393000
1!
1%
1+
#394000
0!
0%
0+
#395000
1!
1%
1+
#396000
0!
0%
0+
#397000
1!
1%
1+
#398000
0!
0%
0+
#399000
1!
1%
1+
#400000
0!
0%
0+
#401000
1!
1%
1+
#402000
0!
0%
0+
#403000
1!
1%
1+
#404000
0!
0%
0+
#405000
1!
1%
1+
#406000
0!
0%
0+
#407000
1!
1%
1+
#408000
0!
0%
0+
#409000
1!
1%
1+
#410000
0!
0%
0+
#411000
1!
1%
1+
#412000
0!
0%
0+
#413000
1!
1%
1+
#414000
0!
0%
0+
#415000
1!
1%
1+
#416000
0!
0%
0+
#417000
1!
1%
1+
#418000
0!
0%
0+
#419000
1!
1%
1+
#420000
0!
0%
0+
#421000
1!
1%
1+
#422000
0!
0%
0+
#423000
1!
1%
1+
#424000
0!
0%
0+
#425000
1!
1%
1+
#426000
0!
0%
0+
#427000
1!
1%
1+
#428000
0!
0%
0+
#429000
1!
1%
1+
#430000
0!
0%
0+
#431000
1!
1%
1+
#432000
0!
0%
0+
#433000
1!
1%
1+
#434000
0!
0%
0+
#435000
1!
1%
1+
#436000
0!
0%
0+
#437000
1!
1%
1+
#438000
0!
0%
0+
#439000
1!
1%
1+
#440000
0!
0%
0+
#441000
1!
1%
1+
#442000
0!
0%
0+
#443000
1!
1%
1+
#444000
0!
0%
0+
#445000
1!
1%
1+
#446000
0!
0%
0+
#447000
1!
1%
1+
#448000
0!
0%
0+
#449000
1!
1%
1+
#450000
0!
0%
0+
#451000
1!
1%
1+
#452000
0!
0%
0+
#453000
1!
1%
1+
#454000
0!
0%
0+
#455000
1!
1%
1+
#456000
0!
0%
0+
#457000
1!
1%
1+
#458000
0!
0%
0+
#459000
1!
1%
1+
#460000
0!
0%
0+
#461000
1!
1%
1+
#462000
0!
0%
0+
#463000
1!
1%
1+
#464000
0!
0%
0+
#465000
1!
1%
1+
#466000
0!
0%
0+
#467000
1!
1%
1+
#468000
0!
0%
0+
#469000
1!
1%
1+
#470000
0!
0%
0+
#471000
1!
1%
1+
#472000
0!
0%
0+
#473000
1!
1%
1+
#474000
0!
0%
0+
#475000
1!
1%
1+
#476000
0!
0%
0+
#477000
1!
1%
1+
#478000
0!
0%
0+
#479000
1!
1%
1+
#480000
0!
0%
0+
#481000
1!
1%
1+
#482000
0!
0%
0+
#483000
1!
1%
1+
#484000
0!
0%
0+
#485000
1!
1%
1+
#486000
0!
0%
0+
#487000
1!
1%
1+
#488000
0!
0%
0+
#489000
1!
1%
1+
#490000
0!
0%
0+
#491000
1!
1%
1+
#492000
0!
0%
0+
#493000
1!
1%
1+
#494000
0!
0%
0+
#495000
1!
1%
1+
#496000
0!
0%
0+
#497000
1!
1%
1+
#498000
0!
0%
0+
#499000
1!
1%
1+
#500000
0!
0%
0+
#501000
1!
1%
1+
#502000
0!
0%
0+
#503000
1!
1%
1+
#504000
0!
0%
0+
#505000
1!
1%
1+
#506000
0!
0%
0+
#507000
1!
1%
1+
#508000
0!
0%
0+
#509000
1!
1%
1+
#510000
0!
0%
0+
#511000
1!
1%
1+
#512000
0!
0%
0+
#513000
1!
1%
1+
#514000
0!
0%
0+
#515000
1!
1%
1+
#516000
0!
0%
0+
#517000
1!
1%
1+
#518000
0!
0%
0+
#519000
1!
1%
1+
#520000
0!
0%
0+
#521000
1!
1%
1+
#522000
0!
0%
0+
#523000
1!
1%
1+
#524000
0!
0%
0+
#525000
1!
1%
1+
#526000
0!
0%
0+
#527000
1!
1%
1+
#528000
0!
0%
0+
#529000
1!
1%
1+
#530000
0!
0%
0+
#531000
1!
1%
1+
#532000
0!
0%
0+
#533000
1!
1%
1+
#534000
0!
0%
0+
#535000
1!
1%
1+
#536000
0!
0%
0+
#537000
1!
1%
1+
#538000
0!
0%
0+
#539000
1!
1%
1+
#540000
0!
0%
0+
#541000
1!
1%
1+
#542000
0!
0%
0+
#543000
1!
1%
1+
#544000
0!
0%
0+
#545000
1!
1%
1+
#546000
0!
0%
0+
#547000
1!
1%
1+
#548000
0!
0%
0+
#549000
1!
1%
1+
#550000
0!
0%
0+
#551000
1!
1%
1+
#552000
0!
0%
0+
#553000
1!
1%
1+
#554000
0!
0%
0+
#555000
1!
1%
1+
#556000
0!
0%
0+
#557000
1!
1%
1+
#558000
0!
0%
0+
#559000
1!
1%
1+
#560000
0!
0%
0+
#561000
1!
1%
1+
#562000
0!
0%
0+
#563000
1!
1%
1+
#564000
0!
0%
0+
#565000
1!
1%
1+
#566000
0!
0%
0+
#567000
1!
1%
1+
#568000
0!
0%
0+
#569000
1!
1%
1+
#570000
0!
0%
0+
#571000
1!
1%
1+
#572000
0!
0%
0+
#573000
1!
1%
1+
#574000
0!
0%
0+
#575000
1!
1%
1+
#576000
0!
0%
0+
#577000
1!
1%
1+
#578000
0!
0%
0+
#579000
1!
1%
1+
#580000
0!
0%
0+
#581000
1!
1%
1+
#582000
0!
0%
0+
#583000
1!
1%
1+
#584000
0!
0%
0+
#585000
1!
1%
1+
#586000
0!
0%
0+
#587000
1!
1%
1+
#588000
0!
0%
0+
#589000
1!
1%
1+
#590000
0!
0%
0+
#591000
1!
1%
1+
#592000
0!
0%
0+
#593000
1!
1%
1+
#594000
0!
0%
0+
#595000
1!
1%
1+
#596000
0!
0%
0+
#597000
1!
1%
1+
#598000
0!
0%
0+
#599000
1!
1%
1+
#600000
0!
0%
0+
#601000
1!
1%
1+
#602000
0!
0%
0+
#603000
1!
1%
1+
#604000
0!
0%
0+
#605000
1!
1%
1+
#606000
0!
0%
0+
#607000
1!
1%
1+
#608000
0!
0%
0+
#609000
1!
1%
1+
#610000
0!
0%
0+
#611000
1!
1%
1+
#612000
0!
0%
0+
#613000
1!
1%
1+
#614000
0!
0%
0+
#615000
1!
1%
1+
#616000
0!
0%
0+
#617000
1!
1%
1+
#618000
0!
0%
0+
#619000
1!
1%
1+
#620000
0!
0%
0+
#621000
1!
1%
1+
#622000
0!
0%
0+
#623000
1!
1%
1+
#624000
0!
0%
0+
#625000
1!
1%
1+
#626000
0!
0%
0+
#627000
1!
1%
1+
#628000
0!
0%
0+
#629000
1!
1%
1+
#630000
0!
0%
0+
#631000
1!
1%
1+
#632000
0!
0%
0+
#633000
1!
1%
1+
#634000
0!
0%
0+
#635000
1!
1%
1+
#636000
0!
0%
0+
#637000
1!
1%
1+
#638000
0!
0%
0+
#639000
1!
1%
1+
#640000
0!
0%
0+
#641000
1!
1%
1+
#642000
0!
0%
0+
#643000
1!
1%
1+
#644000
0!
0%
0+
#645000
1!
1%
1+
#646000
0!
0%
0+
#647000
1!
1%
1+
#648000
0!
0%
0+
#649000
1!
1%
1+
#650000
0!
0%
0+
#651000
1!
1%
1+
#652000
0!
0%
0+
#653000
1!
1%
1+
#654000
0!
0%
0+
#655000
1!
1%
1+
#656000
0!
0%
0+
#657000
1!
1%
1+
#658000
0!
0%
0+
#659000
1!
1%
1+
#660000
0!
0%
0+
#661000
1!
1%
1+
#662000
0!
0%
0+
#663000
1!
1%
1+
#664000
0!
0%
0+
#665000
1!
1%
1+
#666000
0!
0%
0+
#667000
1!
1%
1+
#668000
0!
0%
0+
#669000
1!
1%
1+
#670000
0!
0%
0+
#671000
1!
1%
1+
#672000
0!
0%
0+
#673000
1!
1%
1+
#674000
0!
0%
0+
#675000
1!
1%
1+
#676000
0!
0%
0+
#677000
1!
1%
1+
#678000
0!
0%
0+
#679000
1!
1%
1+
#680000
0!
0%
0+
#681000
1!
1%
1+
#682000
0!
0%
0+
#683000
1!
1%
1+
#684000
0!
0%
0+
#685000
1!
1%
1+
#686000
0!
0%
0+
#687000
1!
1%
1+
#688000
0!
0%
0+
#689000
1!
1%
1+
#690000
0!
0%
0+
#691000
1!
1%
1+
#692000
0!
0%
0+
#693000
1!
1%
1+
#694000
0!
0%
0+
#695000
1!
1%
1+
#696000
0!
0%
0+
#697000
1!
1%
1+
#698000
0!
0%
0+
#699000
1!
1%
1+
#700000
0!
0%
0+
#701000
1!
1%
1+
#702000
0!
0%
0+
#703000
1!
1%
1+
#704000
0!
0%
0+
#705000
1!
1%
1+
#706000
0!
0%
0+
#707000
1!
1%
1+
#708000
0!
0%
0+
#709000
1!
1%
1+
#710000
0!
0%
0+
#711000
1!
1%
1+
#712000
0!
0%
0+
#713000
1!
1%
1+
#714000
0!
0%
0+
#715000
1!
1%
1+
#716000
0!
0%
0+
#717000
1!
1%
1+
#718000
0!
0%
0+
#719000
1!
1%
1+
#720000
0!
0%
0+
#721000
1!
1%
1+
#722000
0!
0%
0+
#723000
1!
1%
1+
#724000
0!
0%
0+
#725000
1!
1%
1+
#726000
0!
0%
0+
#727000
1!
1%
1+
#728000
0!
0%
0+
#729000
1!
1%
1+
#730000
0!
0%
0+
#731000
1!
1%
1+
#732000
0!
0%
0+
#733000
1!
1%
1+
#734000
0!
0%
0+
#735000
1!
1%
1+
#736000
0!
0%
0+
#737000
1!
1%
1+
#738000
0!
0%
0+
#739000
1!
1%
1+
#740000
0!
0%
0+
#741000
1!
1%
1+
#742000
0!
0%
0+
#743000
1!
1%
1+
#744000
0!
0%
0+
#745000
1!
1%
1+
#746000
0!
0%
0+
#747000
1!
1%
1+
#748000
0!
0%
0+
#749000
1!
1%
1+
#750000
0!
0%
0+
#751000
1!
1%
1+
#752000
0!
0%
0+
#753000
1!
1%
1+
#754000
0!
0%
0+
#755000
1!
1%
1+
#756000
0!
0%
0+
#757000
1!
1%
1+
#758000
0!
0%
0+
#759000
1!
1%
1+
#760000
0!
0%
0+
#761000
1!
1%
1+
#762000
0!
0%
0+
#763000
1!
1%
1+
#764000
0!
0%
0+
#765000
1!
1%
1+
#766000
0!
0%
0+
#767000
1!
1%
1+
#768000
0!
0%
0+
#769000
1!
1%
1+
#770000
0!
0%
0+
#771000
1!
1%
1+
#772000
0!
0%
0+
#773000
1!
1%
1+
#774000
0!
0%
0+
#775000
1!
1%
1+
#776000
0!
0%
0+
#777000
1!
1%
1+
#778000
0!
0%
0+
#779000
1!
1%
1+
#780000
0!
0%
0+
#781000
1!
1%
1+
#782000
0!
0%
0+
#783000
1!
1%
1+
#784000
0!
0%
0+
#785000
1!
1%
1+
#786000
0!
0%
0+
#787000
1!
1%
1+
#788000
0!
0%
0+
#789000
1!
1%
1+
#790000
0!
0%
0+
#791000
1!
1%
1+
#792000
0!
0%
0+
#793000
1!
1%
1+
#794000
0!
0%
0+
#795000
1!
1%
1+
#796000
0!
0%
0+
#797000
1!
1%
1+
#798000
0!
0%
0+
#799000
1!
1%
1+
#800000
0!
0%
0+
#801000
1!
1%
1+
#802000
0!
0%
0+
#803000
1!
1%
1+
#804000
0!
0%
0+
#805000
1!
1%
1+
#806000
0!
0%
0+
#807000
1!
1%
1+
#808000
0!
0%
0+
#809000
1!
1%
1+
#810000
0!
0%
0+
#811000
1!
1%
1+
#812000
0!
0%
0+
#813000
1!
1%
1+
#814000
0!
0%
0+
#815000
1!
1%
1+
#816000
0!
0%
0+
#817000
1!
1%
1+
#818000
0!
0%
0+
#819000
1!
1%
1+
#820000
0!
0%
0+
#821000
1!
1%
1+
#822000
0!
0%
0+
#823000
1!
1%
1+
#824000
0!
0%
0+
#825000
1!
1%
1+
#826000
0!
0%
0+
#827000
1!
1%
1+
#828000
0!
0%
0+
#829000
1!
1%
1+
#830000
0!
0%
0+
#831000
1!
1%
1+
#832000
0!
0%
0+
#833000
1!
1%
1+
#834000
0!
0%
0+
#835000
1!
1%
1+
#836000
0!
0%
0+
#837000
1!
1%
1+
#838000
0!
0%
0+
#839000
1!
1%
1+
#840000
0!
0%
0+
#841000
1!
1%
1+
#842000
0!
0%
0+
#843000
1!
1%
1+
#844000
0!
0%
0+
#845000
1!
1%
1+
#846000
0!
0%
0+
#847000
1!
1%
1+
#848000
0!
0%
0+
#849000
1!
1%
1+
#850000
0!
0%
0+
#851000
1!
1%
1+
#852000
0!
0%
0+
#853000
1!
1%
1+
#854000
0!
0%
0+
#855000
1!
1%
1+
#856000
0!
0%
0+
#857000
1!
1%
1+
#858000
0!
0%
0+
#859000
1!
1%
1+
#860000
0!
0%
0+
#861000
1!
1%
1+
#862000
0!
0%
0+
#863000
1!
1%
1+
#864000
0!
0%
0+
#865000
1!
1%
1+
#866000
0!
0%
0+
#867000
1!
1%
1+
#868000
0!
0%
0+
#869000
1!
1%
1+
#870000
0!
0%
0+
#871000
1!
1%
1+
#872000
0!
0%
0+
#873000
1!
1%
1+
#874000
0!
0%
0+
#875000
1!
1%
1+
#876000
0!
0%
0+
#877000
1!
1%
1+
#878000
0!
0%
0+
#879000
1!
1%
1+
#880000
0!
0%
0+
#881000
1!
1%
1+
#882000
0!
0%
0+
#883000
1!
1%
1+
#884000
0!
0%
0+
#885000
1!
1%
1+
#886000
0!
0%
0+
#887000
1!
1%
1+
#888000
0!
0%
0+
#889000
1!
1%
1+
#890000
0!
0%
0+
#891000
1!
1%
1+
#892000
0!
0%
0+
#893000
1!
1%
1+
#894000
0!
0%
0+
#895000
1!
1%
1+
#896000
0!
0%
0+
#897000
1!
1%
1+
#898000
0!
0%
0+
#899000
1!
1%
1+
#900000
0!
0%
0+
#901000
1!
1%
1+
#902000
0!
0%
0+
#903000
1!
1%
1+
#904000
0!
0%
0+
#905000
1!
1%
1+
#906000
0!
0%
0+
#907000
1!
1%
1+
#908000
0!
0%
0+
#909000
1!
1%
1+
#910000
0!
0%
0+
#911000
1!
1%
1+
#912000
0!
0%
0+
#913000
1!
1%
1+
#914000
0!
0%
0+
#915000
1!
1%
1+
#916000
0!
0%
0+
#917000
1!
1%
1+
#918000
0!
0%
0+
#919000
1!
1%
1+
#920000
0!
0%
0+
#921000
1!
1%
1+
#922000
0!
0%
0+
#923000
1!
1%
1+
#924000
0!
0%
0+
#925000
1!
1%
1+
#926000
0!
0%
0+
#927000
1!
1%
1+
#928000
0!
0%
0+
#929000
1!
1%
1+
#930000
0!
0%
0+
#931000
1!
1%
1+
#932000
0!
0%
0+
#933000
1!
1%
1+
#934000
0!
0%
0+
#935000
1!
1%
1+
#936000
0!
0%
0+
#937000
1!
1%
1+
#938000
0!
0%
0+
#939000
1!
1%
1+
#940000
0!
0%
0+
#941000
1!
1%
1+
#942000
0!
0%
0+
#943000
1!
1%
1+
#944000
0!
0%
0+
#945000
1!
1%
1+
#946000
0!
0%
0+
#947000
1!
1%
1+
#948000
0!
0%
0+
#949000
1!
1%
1+
#950000
0!
0%
0+
#951000
1!
1%
1+
#952000
0!
0%
0+
#953000
1!
1%
1+
#954000
0!
0%
0+
#955000
1!
1%
1+
#956000
0!
0%
0+
#957000
1!
1%
1+
#958000
0!
0%
0+
#959000
1!
1%
1+
#960000
0!
0%
0+
#961000
1!
1%
1+
#962000
0!
0%
0+
#963000
1!
1%
1+
#964000
0!
0%
0+
#965000
1!
1%
1+
#966000
0!
0%
0+
#967000
1!
1%
1+
#968000
0!
0%
0+
#969000
1!
1%
1+
#970000
0!
0%
0+
#971000
1!
1%
1+
#972000
0!
0%
0+
#973000
1!
1%
1+
#974000
0!
0%
0+
#975000
1!
1%
1+
#976000
0!
0%
0+
#977000
1!
1%
1+
#978000
0!
0%
0+
#979000
1!
1%
1+
#980000
0!
0%
0+
#981000
1!
1%
1+
#982000
0!
0%
0+
#983000
1!
1%
1+
#984000
0!
0%
0+
#985000
1!
1%
1+
#986000
0!
0%
0+
#987000
1!
1%
1+
#988000
0!
0%
0+
#989000
1!
1%
1+
#990000
0!
0%
0+
#991000
1!
1%
1+
#992000
0!
0%
0+
#993000
1!
1%
1+
#994000
0!
0%
0+
#995000
1!
1%
1+
#996000
0!
0%
0+
#997000
1!
1%
1+
#998000
0!
0%
0+
#999000
1!
1%
1+
#1000000
0!
0%
0+
